library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity pompa is
    port (
        signal clk : in std_logic;
        
    );
end entity pompa;

architecture rtl of pompa is
    
begin
    
    
    
end architecture rtl;